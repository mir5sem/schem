`timescale 1ns / 1ps

/*
???  ??1  ??2  ???

??????? MUL: 4 ??? 4 ??? 4 ??? 4 ???
XNOR: 4 ??? 4 ??? 4 ??? 4 ???

??? ????????? ????????? 
MOV: 4 ??? 4 ??? 4 ???

JUMP: ??? 0000 (8 ??? ????? ???? ??????????)

LOAD: ??? ????? ??? ?????? (4 ???), ??????? (8 ???)
*/

module cpu (
    input clk,
    input reset
);

    parameter DATA_WIDTH = 8; // ??????????? ??????
    parameter ADDR_WIDTH = 8; // ??????????? ??????
    parameter REG_NUM = 16; // ?????????? ?????????
    parameter REG_ADDR_WIDTH = $clog2(REG_NUM); // ??????????? ?????? ?????????
    parameter CMD_WIDTH = 16; // ??????????? ???????

    parameter MUL = 4'b0001; // ?????????
    parameter XNOR = 4'b0010; // ????????? ???????????????
    parameter MOVE = 4'b0011; // ??????????? ?? ???????? ??? ? ??????? ???
    parameter JUMP = 4'b0100; // ???????? ???????
    parameter LOAD = 4'b0101; // ???????? ???????? ? ?????? ??????

    reg [DATA_WIDTH-1:0] data_memory[0:255];
    reg [CMD_WIDTH-1:0] mem_cmd[0:255];

    reg [ADDR_WIDTH-1:0] pc;
    reg [CMD_WIDTH-1:0] cmd_reg;

    wire [DATA_WIDTH-1:0] operand1, operand2;
    reg [DATA_WIDTH-1:0] result;

    reg wen;
    reg [REG_ADDR_WIDTH-1:0] reg_addr_write, reg_addr1, reg_addr2;
    reg [DATA_WIDTH-1:0] reg_data_in;
    wire [DATA_WIDTH-1:0] reg_operand1, reg_operand2;

    reg_file #(.DATA_WIDTH(DATA_WIDTH), .REG_FILE_SIZE(REG_NUM), .ADDR_WIDTH(REG_ADDR_WIDTH)) reg1 (
        .clk(clk), .reset(reset), .wen(wen), .data_in(reg_data_in), .addr_write(reg_addr_write), .addr_a(reg_addr1), .addr_b(reg_addr2), .operand_a(reg_operand1), .operand_b(reg_operand2));

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            pc <= 0;
        end else begin
            // ?????? 0
            cmd_reg <= mem_cmd[pc];
            pc <= pc + 1;

            // ?????? 1
            case (cmd_reg[15:12])
                MUL: begin
                    // ?????????: operand1 * operand2 -> result
                    reg_addr1 <= cmd_reg[11:8];
                    reg_addr2 <= cmd_reg[7:4];
                    reg_addr_write <= cmd_reg[3:0];
                    wen <= 1;
                    reg_data_in <= reg_operand1 * reg_operand2;
                end
                XNOR: begin
                    // ????????? ???????????????: ~(operand1 ^ operand2) -> result
                    reg_addr1 <= cmd_reg[11:8];
                    reg_addr2 <= cmd_reg[7:4];
                    reg_addr_write <= cmd_reg[3:0];
                    wen <= 1;
                    reg_data_in <= ~(reg_operand1 ^ reg_operand2);
                end
                MOVE: begin
                    // ??????????? ???????? ?? ?????? ???????? ? ??????
                    reg_addr1 <= cmd_reg[7:4];
                    reg_addr_write <= cmd_reg[11:8];
                    wen <= 1;
                    reg_data_in <= reg_operand1;
                end
                JUMP: begin
                    // ???????? ???????
                    if (result > 0) begin
                        pc <= cmd_reg[7:0];
                    end
                end
                LOAD: begin
                    // ???????? ???????? ? ?????? ??????
                    data_memory[cmd_reg[11:8]] <= cmd_reg[7:0];
                end
                default: begin
                    // ?? ?????????
                    wen <= 0;
                    reg_addr1 <= cmd_reg[11:8];
                    reg_addr2 <= cmd_reg[7:4];
                    reg_addr_write <= cmd_reg[3:0];
                    reg_data_in <= reg_operand1 * reg_operand2;
                end
            endcase
        end
    end

endmodule
