assign cos_table[00] = 16'b1000000000000000;
assign cos_table[01] = 16'b0111111111011000;
assign cos_table[02] = 16'b0111111101100010;
assign cos_table[03] = 16'b0111111010011101;
assign cos_table[04] = 16'b0111110110001010;
assign cos_table[05] = 16'b0111110000101001;
assign cos_table[06] = 16'b0111101001111101;
assign cos_table[07] = 16'b0111100010000100;
assign cos_table[08] = 16'b0111011001000001;
assign cos_table[09] = 16'b0111001110110101;
assign cos_table[10] = 16'b0111000011100010;
assign cos_table[11] = 16'b0110110111001010;
assign cos_table[12] = 16'b0110101001101101;
assign cos_table[13] = 16'b0110011011001111;
assign cos_table[14] = 16'b0110001011110010;
assign cos_table[15] = 16'b0101111011010111;
assign cos_table[16] = 16'b0101101010000010;
assign cos_table[17] = 16'b0101010111110101;
assign cos_table[18] = 16'b0101000100110011;
assign cos_table[19] = 16'b0100110000111111;
assign cos_table[20] = 16'b0100011100011100;
assign cos_table[21] = 16'b0100000111001110;
assign cos_table[22] = 16'b0011110001010110;
assign cos_table[23] = 16'b0011011010111010;
assign cos_table[24] = 16'b0011000011111011;
assign cos_table[25] = 16'b0010101100011111;
assign cos_table[26] = 16'b0010010100101000;
assign cos_table[27] = 16'b0001111100011001;
assign cos_table[28] = 16'b0001100011111000;
assign cos_table[29] = 16'b0001001011001000;
assign cos_table[30] = 16'b0000110010001011;
assign cos_table[31] = 16'b0000011001000111;
assign cos_table[32] = 16'b0000000000000000;
assign cos_table[33] = 16'b0000011001000111;
assign cos_table[34] = 16'b0000110010001011;
assign cos_table[35] = 16'b0001001011001000;
assign cos_table[36] = 16'b0001100011111000;
assign cos_table[37] = 16'b0001111100011001;
assign cos_table[38] = 16'b0010010100101000;
assign cos_table[39] = 16'b0010101100011111;
assign cos_table[40] = 16'b0011000011111011;
assign cos_table[41] = 16'b0011011010111010;
assign cos_table[42] = 16'b0011110001010110;
assign cos_table[43] = 16'b0100000111001110;
assign cos_table[44] = 16'b0100011100011100;
assign cos_table[45] = 16'b0100110000111111;
assign cos_table[46] = 16'b0101000100110011;
assign cos_table[47] = 16'b0101010111110101;
assign cos_table[48] = 16'b0101101010000010;
assign cos_table[49] = 16'b0101111011010111;
assign cos_table[50] = 16'b0110001011110010;
assign cos_table[51] = 16'b0110011011001111;
assign cos_table[52] = 16'b0110101001101101;
assign cos_table[53] = 16'b0110110111001010;
assign cos_table[54] = 16'b0111000011100010;
assign cos_table[55] = 16'b0111001110110101;
assign cos_table[56] = 16'b0111011001000001;
assign cos_table[57] = 16'b0111100010000100;
assign cos_table[58] = 16'b0111101001111101;
assign cos_table[59] = 16'b0111110000101001;
assign cos_table[60] = 16'b0111110110001010;
assign cos_table[61] = 16'b0111111010011101;
assign cos_table[62] = 16'b0111111101100010;
assign cos_table[63] = 16'b0111111111011000;
assign cos_table[64] = 16'b1000000000000000;
assign cos_table[65] = 16'b0111111111011000;
assign cos_table[66] = 16'b0111111101100010;
assign cos_table[67] = 16'b0111111010011101;
assign cos_table[68] = 16'b0111110110001010;
assign cos_table[69] = 16'b0111110000101001;
assign cos_table[70] = 16'b0111101001111101;
assign cos_table[71] = 16'b0111100010000100;
assign cos_table[72] = 16'b0111011001000001;
assign cos_table[73] = 16'b0111001110110101;
assign cos_table[74] = 16'b0111000011100010;
assign cos_table[75] = 16'b0110110111001010;
assign cos_table[76] = 16'b0110101001101101;
assign cos_table[77] = 16'b0110011011001111;
assign cos_table[78] = 16'b0110001011110010;
assign cos_table[79] = 16'b0101111011010111;
assign cos_table[80] = 16'b0101101010000010;
assign cos_table[81] = 16'b0101010111110101;
assign cos_table[82] = 16'b0101000100110011;
assign cos_table[83] = 16'b0100110000111111;
assign cos_table[84] = 16'b0100011100011100;
assign cos_table[85] = 16'b0100000111001110;
assign cos_table[86] = 16'b0011110001010110;
assign cos_table[87] = 16'b0011011010111010;
assign cos_table[88] = 16'b0011000011111011;
assign cos_table[89] = 16'b0010101100011111;
assign cos_table[90] = 16'b0010010100101000;
assign cos_table[91] = 16'b0001111100011001;
assign cos_table[92] = 16'b0001100011111000;
assign cos_table[93] = 16'b0001001011001000;
assign cos_table[94] = 16'b0000110010001011;
assign cos_table[95] = 16'b0000011001000111;
assign cos_table[96] = 16'b0000000000000000;
assign cos_table[97] = 16'b0000011001000111;
assign cos_table[98] = 16'b0000110010001011;
assign cos_table[99] = 16'b0001001011001000;
assign cos_table[100] = 16'b0001100011111000;
assign cos_table[101] = 16'b0001111100011001;
assign cos_table[102] = 16'b0010010100101000;
assign cos_table[103] = 16'b0010101100011111;
assign cos_table[104] = 16'b0011000011111011;
assign cos_table[105] = 16'b0011011010111010;
assign cos_table[106] = 16'b0011110001010110;
assign cos_table[107] = 16'b0100000111001110;
assign cos_table[108] = 16'b0100011100011100;
assign cos_table[109] = 16'b0100110000111111;
assign cos_table[110] = 16'b0101000100110011;
assign cos_table[111] = 16'b0101010111110101;
assign cos_table[112] = 16'b0101101010000010;
assign cos_table[113] = 16'b0101111011010111;
assign cos_table[114] = 16'b0110001011110010;
assign cos_table[115] = 16'b0110011011001111;
assign cos_table[116] = 16'b0110101001101101;
assign cos_table[117] = 16'b0110110111001010;
assign cos_table[118] = 16'b0111000011100010;
assign cos_table[119] = 16'b0111001110110101;
assign cos_table[120] = 16'b0111011001000001;
assign cos_table[121] = 16'b0111100010000100;
assign cos_table[122] = 16'b0111101001111101;
assign cos_table[123] = 16'b0111110000101001;
assign cos_table[124] = 16'b0111110110001010;
assign cos_table[125] = 16'b0111111010011101;
assign cos_table[126] = 16'b0111111101100010;
assign cos_table[127] = 16'b0111111111011000;
